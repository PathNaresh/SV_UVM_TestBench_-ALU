interface my_interface(input logic clock);

  logic reset;
  logic [2:0] a, b;
  logic sel;
  logic [3:0] result;

endinterface
